module datapath();
    
endmodule