// `define INPUT_IMAGES 
// ``define  Fill_value
