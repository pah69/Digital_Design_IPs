//  Package: ALU_pkg
//
package ALU_pkg;
    //  Group: Typedefs
    typedef enum {
        Add,
        Sub,
        LeftShift,
        RightShiftArith,
        RightShiftLogic,
        And,
        Or,
        Xor,
        Equal
      } OpCode;

    //  Group: Parameters
    

    
endpackage: ALU_pkg
