module pc_mux (
    input logic pc_src,
    input logic [31:0] pc
)
endmodule