//  Package: pkg
//
package alu_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  //  Group: Typedefs
  `include "seq_item.svh"
  `include "base_seq.svh"
  `include "sequencer.svh"
  `include "driver.svh"
  `include "monitor.svh"
  `include "scoreboard.svh"
  `include "agent.svh"
  `include "env.svh"
  `include "base_test.sv"
  //  Group: Parameters



endpackage
