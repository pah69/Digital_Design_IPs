module FIFO #(
    parameter  DataWidth = 32,
    parameter  Depth     = 8,
    localparam PtrWidth  = $clog2(Depth)
  ) (
    input  logic                 clk,
    input  logic                 rstN,
    input  logic                 writeEn,
    input  logic [DataWidth-1:0] writeData,
    input  logic                 readEn,
    output logic [DataWidth-1:0] readData,
    output logic                 full,
    output logic                 empty
  );
  
    logic [DataWidth-1:0] mem[Depth];
    logic [PtrWidth:0] wrPtr, wrPtrNext;
    logic [PtrWidth:0] rdPtr, rdPtrNext;
  
    always_comb begin
      wrPtrNext = wrPtr;
      rdPtrNext = rdPtr;
      if (writeEn) begin
        wrPtrNext = wrPtr + 1;
      end
      if (readEn) begin
        rdPtrNext = rdPtr + 1;
      end
    end
  
    always_ff @(posedge clk or negedge rstN) begin
      if (!rstN) begin
        wrPtr <= '0;
        rdPtr <= '0;
      end else begin
        wrPtr <= wrPtrNext;
        rdPtr <= rdPtrNext;
      end
  
      mem[wrPtr[PtrWidth-1:0]] <= writeData;
    end
  
    assign readData = mem[rdPtr[PtrWidth-1:0]];
  
    assign empty = (wrPtr[PtrWidth] == rdPtr[PtrWidth]) && (wrPtr[PtrWidth-1:0] == rdPtr[PtrWidth-1:0]);
    assign full  = (wrPtr[PtrWidth] != rdPtr[PtrWidth]) && (wrPtr[PtrWidth-1:0] == rdPtr[PtrWidth-1:0]);
  
  endmodule