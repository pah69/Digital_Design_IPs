
// Up or Down Counter

