
// Modulo Counter
