module controller();



    main_decoder();

    alu_decoder();

    

endmodule