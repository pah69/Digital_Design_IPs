module input_layer#(

) (
    input 
)
