module test(
    port_list
);
    
endmodule