module imm_gen(
    input logic [31:0] instruction,
    output 
);
    
endmodule