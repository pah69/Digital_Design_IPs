module FIFO(
    input logic a;
    output logic out;
);
    
endmodule